module BK0717A();
endmodule